module vga_graphics(
    input  wire [9:0] x,
    input  wire [9:0] y,
    input  wire en,
    output reg [3:0] red,
    output reg [3:0] green,
    output reg [3:0] blue
);

localparam Wide = 213;   // 640 / 3
localparam High = 160;   // 480 / 3
localparam LINE_W =   5;

    wire [9:0] rel_x = x % Wide;
    wire [9:0] rel_y = y % High;

wire border =
       (rel_x < LINE_W)
    || (rel_x >= Wide - LINE_W)
    || (rel_y < LINE_W)
    || (rel_y >= High - LINE_W);

always @(*) begin
    if (!en) begin // black
        red   = 4'h0;
        green = 4'h0;
        blue  = 4'h0;
    end else if (border) begin //black
        red   = 4'h0;
        green = 4'h0;
        blue  = 4'h0;
    end else begin // white
        red   = 4'hF;
        green = 4'hF;
        blue  = 4'hF;
    end
end

endmodule



