module clk25_chain (
    input  wire clk,
    input  wire reset,
    output wire clk25
);
    wire q0;

    counter #(
        .MaxCount  (1),
        .DataWidth (1)
    ) U_DIV2_1 (
        .clk   (clk),
        .reset (reset),
        .en    (1'b1),
        .Q     (q0),
        .TC    ()
    );

    counter #(
        .MaxCount  (1),
        .DataWidth (1)
    ) U_DIV2_2 (
        .clk   (clk),
        .reset (reset),
        .en    (q0),
        .Q     (clk25),
        .TC    ()
    );

endmodule
