module uart_controller (
    input  wire       clk,
    input  wire       reset,
    input  wire       rx_in,
    output wire       up,
    output wire       down,
    output wire       left,
    output wire       right,
    output wire       enter,
    output wire       space
);

    wire [7:0] rx_data;
    wire rx_valid;

    uart_rx u_rx (
        .clk(clk),
        .reset(reset),
        .rx_in(rx_in),
        .rx_out(rx_data),
        .rx_valid(rx_valid)
    );

    key_decoder u_decoder (
        .clk(clk),
        .reset(reset),
        .data(rx_data),
        .rx_valid(rx_valid),
        .up(up),
        .down(down),
        .left(left),
        .right(right),
        .enter(enter),
        .space(space)
    );

endmodule