
module vga_top (
    input  wire       clk25,          // 25MHz clock from external source
    input  wire       reset,
    input  wire [17:0] sw, // Use 18-bit input for 9 cells (2 bits each)
    input  wire [8:0] cell_select_flag, // One-hot encoding for cursor position
    output wire       VGA_HS,
    output wire       VGA_VS,
    output wire [3:0] VGA_R,
    output wire [3:0] VGA_G,
    output wire [3:0] VGA_B
);

    // VGA sync signals and coordinates
    wire [9:0] x;
    wire [9:0] y;
    wire       en;
    vga_sync u_sync (
        .clk      (clk25),
        .reset    (reset), // Use the main reset directly
        .x        (x),
        .y        (y),
        .hsync    (VGA_HS),
        .vsync    (VGA_VS),
        .en       (en)
    );

    // Graphics generator
    vga_graphics u_grp (
        .clk      (clk25),
        .reset    (reset), // Use the main reset directly
        .x        (x),
        .y        (y),
        .en       (en),
        .sw       (sw),
        .cell_select_flag (cell_select_flag),
        .red      (VGA_R),
        .green    (VGA_G),
        .blue     (VGA_B)
    );

endmodule
